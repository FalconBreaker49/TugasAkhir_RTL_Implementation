// File Testbench untuk module Reward_Decider

