// File Testbench untuk module Control Unit. 
