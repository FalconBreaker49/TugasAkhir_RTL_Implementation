// File Testbench untuk module Policy Generator (PG). 
